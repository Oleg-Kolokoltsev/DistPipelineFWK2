RC transient process
* Testing transient modelling with an LC contour

* --------- devices ---------
C_C1 0 N_2 1u
R_R2 N_1 N_3 4
L_L1 N_2 N_1 500u
V_V1 N_3 0 DC 0V AC 1 PULSE(-1 1 0 0m 0m 1m 2m)

.TRAN 1e-5 0.500 0 1e-5
.save V(N_2) V(N_3)

.end